`ifndef _base_
`define _base_

class base_pkt;
randc bit Din;
bit rst;
bit Q;
endclass
`endif
